library verilog;
use verilog.vl_types.all;
entity MaquinaEst2_vlg_vec_tst is
end MaquinaEst2_vlg_vec_tst;
