

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;


ENTITY testbench_Restador4Bit is

end testbench_Restador4Bit;

