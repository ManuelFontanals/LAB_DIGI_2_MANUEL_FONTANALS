library verilog;
use verilog.vl_types.all;
entity RestadorCompleto_vlg_check_tst is
    port(
        o_bout          : in     vl_logic;
        o_res           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end RestadorCompleto_vlg_check_tst;
