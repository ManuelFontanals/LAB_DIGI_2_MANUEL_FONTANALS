library verilog;
use verilog.vl_types.all;
entity ConexionMasterSlave_vlg_vec_tst is
end ConexionMasterSlave_vlg_vec_tst;
