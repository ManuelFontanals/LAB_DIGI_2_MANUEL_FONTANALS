library verilog;
use verilog.vl_types.all;
entity SumadorCompletoProcess_vlg_vec_tst is
end SumadorCompletoProcess_vlg_vec_tst;
