library verilog;
use verilog.vl_types.all;
entity RestadorCompleto_vlg_vec_tst is
end RestadorCompleto_vlg_vec_tst;
