-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 06 17:26:51 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MaquinaEstado IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z : OUT STD_LOGIC
    );
END MaquinaEstado;

ARCHITECTURE BEHAVIOR OF MaquinaEstado IS
    TYPE type_fstate IS (A,B,D,C);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            Z <= '0';
        ELSE
            Z <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '1')) THEN
                        reg_fstate <= B;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= A;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    IF ((x = '1')) THEN
                        Z <= '0';
                    ELSIF ((x = '0')) THEN
                        Z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= '0';
                    END IF;
                WHEN B =>
                    IF ((x = '0')) THEN
                        reg_fstate <= A;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;

                    IF ((x = '1')) THEN
                        Z <= '0';
                    ELSIF ((x = '0')) THEN
                        Z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= '0';
                    END IF;
                WHEN D =>
                    IF ((x = '0')) THEN
                        reg_fstate <= A;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D;
                    END IF;

                    IF ((x = '1')) THEN
                        Z <= '0';
                    ELSIF ((x = '0')) THEN
                        Z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= '0';
                    END IF;
                WHEN C =>
                    IF ((x = '0')) THEN
                        reg_fstate <= A;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= C;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    IF ((x = '1')) THEN
                        Z <= '1';
                    ELSIF ((x = '0')) THEN
                        Z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        Z <= '0';
                    END IF;
                WHEN OTHERS => 
                    Z <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
