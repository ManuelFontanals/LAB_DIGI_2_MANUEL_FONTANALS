library verilog;
use verilog.vl_types.all;
entity SumadorDefBloq_vlg_vec_tst is
end SumadorDefBloq_vlg_vec_tst;
