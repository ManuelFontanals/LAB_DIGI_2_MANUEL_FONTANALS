-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 06 19:28:42 2024




   --  ACLARACION:
	
   --   ASUMO QUE LAS ENTRADAS VIENEN DE UN CIRCUITO APARTE, NO SINTETIZO EN ESTA FPGA NI CONTADORES, NI REGISTROS ETC, SOLO LA LÓGICA DE SETEO DEL SLAVE




LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ConexionMasterSlave IS
    PORT (
        reset : IN STD_LOGIC := '0';
        SCL : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        Hab_dir : OUT STD_LOGIC;
        Hab_Data : OUT STD_LOGIC;
        ACK : OUT STD_LOGIC
    );
END ConexionMasterSlave;

ARCHITECTURE BEHAVIOR OF ConexionMasterSlave IS
    TYPE type_fstate IS (Idle,DirCheck,WriteOrRead,WaitConec,SaveData,Start);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (SCL,reg_fstate)
    BEGIN
        IF (SCL='1' AND SCL'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,fin_dir,fin_dato,soy)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Idle;
            Hab_dir <= '0';
            Hab_Data <= '0';
            ACK <= '0';
        ELSE
            Hab_dir <= '0';
            Hab_Data <= '0';
            ACK <= '0';
            CASE fstate IS
                WHEN Idle =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Start;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= Idle;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Idle;
                    END IF;

                    Hab_dir <= '0';

                    Hab_Data <= '0';

                    ACK <= '0';
                WHEN DirCheck =>
                    IF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= WriteOrRead;
                    ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Idle;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= DirCheck;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DirCheck;
                    END IF;

                    Hab_dir <= '1';

                    Hab_Data <= '0';

                    ACK <= '0';
                WHEN WriteOrRead =>
                    reg_fstate <= WaitConec;

                    Hab_dir <= '0';

                    Hab_Data <= '0';

                    ACK <= '0';
                WHEN WaitConec =>
                    reg_fstate <= SaveData;

                    Hab_dir <= '0';

                    Hab_Data <= '0';

                    ACK <= '1';
                WHEN SaveData =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= SaveData;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SaveData;
                    END IF;

                    Hab_dir <= '0';

                    Hab_Data <= '1';

                    ACK <= '0';
                WHEN Start =>
                    reg_fstate <= DirCheck;

                    Hab_dir <= '0';

                    Hab_Data <= '0';

                    ACK <= '0';
                WHEN OTHERS => 
                    Hab_dir <= 'X';
                    Hab_Data <= 'X';
                    ACK <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
