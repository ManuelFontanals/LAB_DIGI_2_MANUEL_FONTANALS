library verilog;
use verilog.vl_types.all;
entity SumadorCompletoProcess_vlg_check_tst is
    port(
        o_cout          : in     vl_logic;
        o_res           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SumadorCompletoProcess_vlg_check_tst;
