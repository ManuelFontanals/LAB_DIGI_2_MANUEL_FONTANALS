library verilog;
use verilog.vl_types.all;
entity Parte_A_vlg_vec_tst is
end Parte_A_vlg_vec_tst;
