library verilog;
use verilog.vl_types.all;
entity SumadorCompleto_vlg_vec_tst is
end SumadorCompleto_vlg_vec_tst;
