library verilog;
use verilog.vl_types.all;
entity MaquinaEstado_vlg_vec_tst is
end MaquinaEstado_vlg_vec_tst;
