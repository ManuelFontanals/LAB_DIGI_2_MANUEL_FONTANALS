library ieee;
use ieee.std_logic;

entity Restador6Bit is
Port 