library verilog;
use verilog.vl_types.all;
entity AgrandoA_vlg_vec_tst is
end AgrandoA_vlg_vec_tst;
