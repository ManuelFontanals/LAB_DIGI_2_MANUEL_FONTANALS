library verilog;
use verilog.vl_types.all;
entity TestStateMach_vlg_vec_tst is
end TestStateMach_vlg_vec_tst;
