library verilog;
use verilog.vl_types.all;
entity MaquinaEstado_vlg_check_tst is
    port(
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MaquinaEstado_vlg_check_tst;
