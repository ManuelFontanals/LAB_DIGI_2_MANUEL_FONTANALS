library verilog;
use verilog.vl_types.all;
entity Parte_A_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Parte_A_vlg_check_tst;
